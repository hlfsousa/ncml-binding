netcdf cami_0000-09-01_64x128_L26_c030918 {
dimensions:
	lat = 64 ;
	lon = 128 ;
	lev = 26 ;
	ilev = 27 ;
	time = UNLIMITED ; // (1 currently)
	chars = 8 ;
variables:
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 9.99999961690316e+35 ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 9.99999961690316e+35 ;
	double lev(lev) ;
		lev:long_name = "hybrid level at midpoints (1000*(A+B))" ;
		lev:units = "level" ;
		lev:positive = "down" ;
		lev:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
		lev:formula_terms = "a: hyam b: hybm p0: P0 ps: PS" ;
		lev:_FillValue = 9.99999961690316e+35 ;
	double ilev(ilev) ;
		ilev:long_name = "hybrid level at interfaces (1000*(A+B))" ;
		ilev:units = "level" ;
		ilev:positive = "down" ;
		ilev:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
		ilev:formula_terms = "a: hyai b: hybi p0: P0 ps: PS" ;
		ilev:_FillValue = 9.99999961690316e+35 ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0000-08-29 00:00:00" ;
		time:calendar = "noleap" ;
		time:_FillValue = 9.99999961690316e+35 ;
	double hyai(ilev) ;
		hyai:long_name = "hybrid A coefficient at layer interfaces" ;
		hyai:_FillValue = 9.99999961690316e+35 ;
	double hybi(ilev) ;
		hybi:long_name = "hybrid B coefficient at layer interfaces" ;
		hybi:_FillValue = 9.99999961690316e+35 ;
	double hyam(lev) ;
		hyam:long_name = "hybrid A coefficient at layer midpoints" ;
		hyam:_FillValue = 9.99999961690316e+35 ;
	double hybm(lev) ;
		hybm:long_name = "hybrid B coefficient at layer midpoints" ;
		hybm:_FillValue = 9.99999961690316e+35 ;
	double gw(lat) ;
		gw:long_name = "gauss weights" ;
		gw:_FillValue = 9.99999961690316e+35 ;
	double P0 ;
		P0:long_name = "reference pressure" ;
		P0:units = "Pa" ;
	char date_written(time, chars) ;
	char time_written(time, chars) ;
	int ntrm ;
		ntrm:long_name = "spectral truncation parameter M" ;
	int ntrn ;
		ntrn:long_name = "spectral truncation parameter N" ;
	int ntrk ;
		ntrk:long_name = "spectral truncation parameter K" ;
	int ndbase ;
		ndbase:long_name = "base day" ;
	int nsbase ;
		nsbase:long_name = "seconds of base day" ;
	int nbdate ;
		nbdate:long_name = "base date (YYYYMMDD)" ;
	int nbsec ;
		nbsec:long_name = "seconds of base date" ;
	int mdt ;
		mdt:long_name = "timestep" ;
		mdt:units = "s" ;
	int ndcur(time) ;
		ndcur:long_name = "current day (from base day)" ;
	int nscur(time) ;
		nscur:long_name = "current seconds of current day" ;
	int date(time) ;
		date:long_name = "current date (YYYYMMDD)" ;
	int datesec(time) ;
		datesec:long_name = "current seconds of current date" ;
	int nsteph(time) ;
		nsteph:long_name = "current timestep" ;
	double U(time, lat, lev, lon) ;
		U:long_name = "Zonal wind" ;
		U:units = "m/s" ;
	double V(time, lat, lev, lon) ;
		V:long_name = "Meridional wind" ;
		V:units = "m/s" ;
	double T(time, lat, lev, lon) ;
		T:long_name = "Temperature" ;
		T:units = "K" ;
	double Q(time, lat, lev, lon) ;
		Q:long_name = "Specific humidity" ;
		Q:units = "kg/kg" ;
	double PS(time, lat, lon) ;
		PS:long_name = "Surface pressure" ;
		PS:units = "Pa" ;
	double PHIS(time, lat, lon) ;
		PHIS:long_name = "surface geopotential" ;
		PHIS:units = "M2/S2" ;
		PHIS:_FillValue = 1.e+36 ;
		PHIS:from_hires = "true" ;
	double SGH(time, lat, lon) ;
		SGH:long_name = "orography standard deviation" ;
		SGH:units = "M" ;
		SGH:_FillValue = 1.e+36 ;
		SGH:from_hires = "true" ;
	double LANDM(time, lat, lon) ;
		LANDM:long_name = "land ocean transition mask: ocean (0), continent (1), transition (0-1)" ;
		LANDM:units = "none" ;
		LANDM:_FillValue = 1.e+36 ;
		LANDM:from_hires = "true" ;
	double PBLH(time, lat, lon) ;
		PBLH:long_name = "PBL height" ;
		PBLH:units = "m" ;
	double TPERT(time, lat, lon) ;
		TPERT:long_name = "Perturbation temperature (eddies in PBL)" ;
		TPERT:units = "K" ;
	double QPERT(time, lat, lon) ;
		QPERT:long_name = "Perturbation specific humidity (eddies in PBL)" ;
		QPERT:units = "kg/kg" ;
	double CLOUD(time, lat, lev, lon) ;
		CLOUD:long_name = "Cloud fraction" ;
		CLOUD:units = "fraction" ;
	double QCWAT(time, lat, lev, lon) ;
	double TCWAT(time, lat, lev, lon) ;
	double LCWAT(time, lat, lev, lon) ;
	double TSICERAD(time, lat, lon) ;
	double TS(time, lat, lon) ;
		TS:long_name = "Surface temperature" ;
		TS:units = "K" ;
	double TSICE(time, lat, lon) ;
		TSICE:long_name = "Ice temperature" ;
		TSICE:units = "K" ;
	double TS1(time, lat, lon) ;
		TS1:long_name = "TS1      subsoil temperature" ;
		TS1:units = "K" ;
	double TS2(time, lat, lon) ;
		TS2:long_name = "TS2      subsoil temperature" ;
		TS2:units = "K" ;
	double TS3(time, lat, lon) ;
		TS3:long_name = "TS3      subsoil temperature" ;
		TS3:units = "K" ;
	double TS4(time, lat, lon) ;
		TS4:long_name = "TS4      subsoil temperature" ;
		TS4:units = "K" ;
	double SNOWHICE(time, lat, lon) ;
		SNOWHICE:long_name = "Water equivalent snow depth" ;
		SNOWHICE:units = "m" ;
	double LANDFRAC(time, lat, lon) ;
		LANDFRAC:long_name = "gridbox land fraction" ;
		LANDFRAC:units = "FRAC" ;
		LANDFRAC:_FillValue = 1.e+36 ;
		LANDFRAC:from_hires = "true" ;
	double TBOT(time, lat, lon) ;
		TBOT:long_name = "Lowest model level temperature" ;
		TBOT:units = "K" ;
	double ICEFRAC(time, lat, lon) ;
		ICEFRAC:long_name = "Fraction of sfc area covered by sea-ice" ;
		ICEFRAC:units = "fraction" ;
	double SICTHK(time, lat, lon) ;
		SICTHK:long_name = "Sea ice thickness" ;
		SICTHK:units = "m" ;
	double TSOCN(time, lat, lon) ;
	double CLDLIQ(time, lat, lev, lon) ;
		CLDLIQ:long_name = "Grid box averaged liquid condensate amount" ;
		CLDLIQ:units = "kg/kg" ;
	double CLDICE(time, lat, lev, lon) ;
		CLDICE:long_name = "Grid box averaged ice condensate amount" ;
		CLDICE:units = "kg/kg" ;
	double LANDM_COSLAT(time, lat, lon) ;
		LANDM_COSLAT:long_name = "land ocean transition mask: ocean (0), continent (1), transition (0-1)" ;
		LANDM_COSLAT:units = "none" ;
		LANDM_COSLAT:_FillValue = 1.e+36 ;
		LANDM_COSLAT:from_hires = "true" ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:logname = "olson" ;
		:host = "bb0001en" ;
		:source = "Interpolated from:/fs/cgd/data0/olson/inputIC/newICeul.cam2.i.0000-09-01-00000.nc::CAM" ;
		:case = "cam2run" ;
		:title = "Interpolated from:/fs/cgd/data0/olson/inputIC/newICeul.cam2.i.0000-09-01-00000.nc::atm ver atm, eul ver v013, case newICeul" ;
		:history = "\n",
    "05/07/03 12:15:34 olson:chinookfe:interpic -t SEP1.T42L26.gaussian.template.nc /fs/cgd/data0/olson/inputIC/newICeul.cam2.i.0000-09-01-00000.nc cami_0000-09-01_64x128_L26_c030507.nc\n",
    "definesurf -t /fs/cgd/csm/inputdata/atm/cam1/hrtopo/topo.nc cami_0000-09-01_64x128_L26_c030507.nc\n",
    "definesurf -t /fs/cgd/csm/inputdata/atm/cam2/hrtopo/topo.nc cami_0000-09-01_64x128_L26_c030507.nc\n",
    "definesurf -t /fs/cgd/csm/inputdata/atm/cam2/hrtopo/topo-usgs-10min.nc cami_0000-09-01_64x128_L26_c030507.nc\n",
    "definesurf -t /fs/cgd/csm/inputdata/atm/cam2/hrtopo/topo10min.merged_c030506.nc cami_0000-09-01_64x128_L26_c030507.nc\n",
    "definesurf -t /fs/cgd/csm/inputdata/atm/cam2/hrtopo/topo10min.merged_c030506.nc -l cami_0000-09-01_64x128_L26_c030624.nc.new" ;
		:make_ross = "true" ;
data:

 lat = -87.8637988392335, -85.0965269883176, -82.3129129478865, 
    -79.5256065726595, -76.7368996803684, -73.9475151539897, 
    -71.1577520115874, -68.3677561083132, -65.5776070108279, 
    -62.7873517989631, -59.9970201084913, -57.2066315276433, 
    -54.4161995260863, -51.6257336749383, -48.8352409662506, 
    -46.0447266311017, -43.254194665351, -40.463648178115, -37.6730896290454, 
    -34.8825209937735, -32.091943881744, -29.3013596217627, -26.510769325211, 
    -23.7201739335347, -20.9295742544895, -18.1389709902393, 
    -15.3483647594915, -12.5577561152307, -9.76714555919551, 
    -6.97653355394858, -4.18592053318916, -1.39530691081949, 
    1.39530691081953, 4.18592053318919, 6.97653355394868, 9.76714555919561, 
    12.5577561152307, 15.3483647594915, 18.1389709902394, 20.9295742544895, 
    23.7201739335347, 26.510769325211, 29.3013596217628, 32.0919438817441, 
    34.8825209937734, 37.6730896290454, 40.4636481781151, 43.254194665351, 
    46.0447266311017, 48.8352409662506, 51.6257336749383, 54.4161995260862, 
    57.2066315276433, 59.9970201084913, 62.7873517989631, 65.5776070108278, 
    68.3677561083132, 71.1577520115871, 73.9475151539896, 76.7368996803683, 
    79.5256065726595, 82.3129129478864, 85.0965269883172, 87.8637988392326 ;

 lon = 0, 2.8125, 5.625, 8.4375, 11.25, 14.0625, 16.875, 19.6875, 22.5, 
    25.3125, 28.125, 30.9375, 33.75, 36.5625, 39.375, 42.1875, 45, 47.8125, 
    50.625, 53.4375, 56.25, 59.0625, 61.875, 64.6875, 67.5, 70.3125, 73.125, 
    75.9375, 78.75, 81.5625, 84.375, 87.1875, 90, 92.8125, 95.625, 98.4375, 
    101.25, 104.0625, 106.875, 109.6875, 112.5, 115.3125, 118.125, 120.9375, 
    123.75, 126.5625, 129.375, 132.1875, 135, 137.8125, 140.625, 143.4375, 
    146.25, 149.0625, 151.875, 154.6875, 157.5, 160.3125, 163.125, 165.9375, 
    168.75, 171.5625, 174.375, 177.1875, 180, 182.8125, 185.625, 188.4375, 
    191.25, 194.0625, 196.875, 199.6875, 202.5, 205.3125, 208.125, 210.9375, 
    213.75, 216.5625, 219.375, 222.1875, 225, 227.8125, 230.625, 233.4375, 
    236.25, 239.0625, 241.875, 244.6875, 247.5, 250.3125, 253.125, 255.9375, 
    258.75, 261.5625, 264.375, 267.1875, 270, 272.8125, 275.625, 278.4375, 
    281.25, 284.0625, 286.875, 289.6875, 292.5, 295.3125, 298.125, 300.9375, 
    303.75, 306.5625, 309.375, 312.1875, 315, 317.8125, 320.625, 323.4375, 
    326.25, 329.0625, 331.875, 334.6875, 337.5, 340.3125, 343.125, 345.9375, 
    348.75, 351.5625, 354.375, 357.1875 ;

 lev = 3.54463800000001, 7.38881350000001, 13.967214, 23.944625, 
    37.2302900000001, 53.1146050000002, 70.0591500000003, 85.4391150000003, 
    100.514695, 118.250335, 139.115395, 163.66207, 192.539935, 226.513265, 
    266.481155, 313.501265000001, 368.817980000002, 433.895225000001, 
    510.455255000002, 600.524200000003, 696.796290000003, 787.702060000003, 
    867.160760000001, 929.648875000002, 970.554830000001, 992.5561 ;

 ilev = 2.19406700000001, 4.89520900000001, 9.882418, 18.05201, 29.83724, 
    44.6233400000002, 61.6058700000002, 78.5124300000004, 92.3658000000002, 
    108.66359, 127.83708, 150.393710000001, 176.93043, 208.149440000001, 
    244.87709, 288.08522, 338.917310000001, 398.718650000002, 469.0718, 
    551.838710000003, 649.209690000002, 744.382890000004, 831.021230000001, 
    903.300290000002, 955.997460000003, 985.1122, 1000 ;

 time = 3 ;
}
